`define BEAM_0_ANTENNA_DELAY_0 1
`define BEAM_0_ANTENNA_DELAY_1 4
`define BEAM_0_ANTENNA_DELAY_2 2
`define BEAM_0_ANTENNA_DELAY_3 0
`define BEAM_0_ANTENNA_DELAY_4 3
`define BEAM_0_ANTENNA_DELAY_5 4
`define BEAM_0_ANTENNA_DELAY_6 2
`define BEAM_0_ANTENNA_DELAY_7 0
`define BEAM_1_ANTENNA_DELAY_0 0
`define BEAM_1_ANTENNA_DELAY_1 5
`define BEAM_1_ANTENNA_DELAY_2 3
`define BEAM_1_ANTENNA_DELAY_3 1
`define BEAM_1_ANTENNA_DELAY_4 2
`define BEAM_1_ANTENNA_DELAY_5 4
`define BEAM_1_ANTENNA_DELAY_6 2
`define BEAM_1_ANTENNA_DELAY_7 0
`define BEAM_2_ANTENNA_DELAY_0 0
`define BEAM_2_ANTENNA_DELAY_1 4
`define BEAM_2_ANTENNA_DELAY_2 2
`define BEAM_2_ANTENNA_DELAY_3 0
`define BEAM_2_ANTENNA_DELAY_4 2
`define BEAM_2_ANTENNA_DELAY_5 5
`define BEAM_2_ANTENNA_DELAY_6 3
`define BEAM_2_ANTENNA_DELAY_7 1
`define BEAM_3_ANTENNA_DELAY_0 0
`define BEAM_3_ANTENNA_DELAY_1 5
`define BEAM_3_ANTENNA_DELAY_2 4
`define BEAM_3_ANTENNA_DELAY_3 2
`define BEAM_3_ANTENNA_DELAY_4 2
`define BEAM_3_ANTENNA_DELAY_5 5
`define BEAM_3_ANTENNA_DELAY_6 4
`define BEAM_3_ANTENNA_DELAY_7 2
`define BEAM_4_ANTENNA_DELAY_0 0
`define BEAM_4_ANTENNA_DELAY_1 7
`define BEAM_4_ANTENNA_DELAY_2 5
`define BEAM_4_ANTENNA_DELAY_3 4
`define BEAM_4_ANTENNA_DELAY_4 2
`define BEAM_4_ANTENNA_DELAY_5 6
`define BEAM_4_ANTENNA_DELAY_6 5
`define BEAM_4_ANTENNA_DELAY_7 3
`define BEAM_5_ANTENNA_DELAY_0 0
`define BEAM_5_ANTENNA_DELAY_1 6
`define BEAM_5_ANTENNA_DELAY_2 5
`define BEAM_5_ANTENNA_DELAY_3 3
`define BEAM_5_ANTENNA_DELAY_4 2
`define BEAM_5_ANTENNA_DELAY_5 7
`define BEAM_5_ANTENNA_DELAY_6 5
`define BEAM_5_ANTENNA_DELAY_7 4
`define BEAM_6_ANTENNA_DELAY_0 0
`define BEAM_6_ANTENNA_DELAY_1 8
`define BEAM_6_ANTENNA_DELAY_2 6
`define BEAM_6_ANTENNA_DELAY_3 5
`define BEAM_6_ANTENNA_DELAY_4 2
`define BEAM_6_ANTENNA_DELAY_5 8
`define BEAM_6_ANTENNA_DELAY_6 6
`define BEAM_6_ANTENNA_DELAY_7 5
`define BEAM_7_ANTENNA_DELAY_0 0
`define BEAM_7_ANTENNA_DELAY_1 8
`define BEAM_7_ANTENNA_DELAY_2 7
`define BEAM_7_ANTENNA_DELAY_3 6
`define BEAM_7_ANTENNA_DELAY_4 1
`define BEAM_7_ANTENNA_DELAY_5 7
`define BEAM_7_ANTENNA_DELAY_6 6
`define BEAM_7_ANTENNA_DELAY_7 5
`define BEAM_8_ANTENNA_DELAY_0 0
`define BEAM_8_ANTENNA_DELAY_1 8
`define BEAM_8_ANTENNA_DELAY_2 7
`define BEAM_8_ANTENNA_DELAY_3 6
`define BEAM_8_ANTENNA_DELAY_4 2
`define BEAM_8_ANTENNA_DELAY_5 9
`define BEAM_8_ANTENNA_DELAY_6 8
`define BEAM_8_ANTENNA_DELAY_7 7
`define BEAM_9_ANTENNA_DELAY_0 0
`define BEAM_9_ANTENNA_DELAY_1 10
`define BEAM_9_ANTENNA_DELAY_2 9
`define BEAM_9_ANTENNA_DELAY_3 8
`define BEAM_9_ANTENNA_DELAY_4 2
`define BEAM_9_ANTENNA_DELAY_5 10
`define BEAM_9_ANTENNA_DELAY_6 9
`define BEAM_9_ANTENNA_DELAY_7 8
`define BEAM_10_ANTENNA_DELAY_0 0
`define BEAM_10_ANTENNA_DELAY_1 10
`define BEAM_10_ANTENNA_DELAY_2 10
`define BEAM_10_ANTENNA_DELAY_3 9
`define BEAM_10_ANTENNA_DELAY_4 1
`define BEAM_10_ANTENNA_DELAY_5 9
`define BEAM_10_ANTENNA_DELAY_6 9
`define BEAM_10_ANTENNA_DELAY_7 8
`define BEAM_11_ANTENNA_DELAY_0 0
`define BEAM_11_ANTENNA_DELAY_1 9
`define BEAM_11_ANTENNA_DELAY_2 9
`define BEAM_11_ANTENNA_DELAY_3 8
`define BEAM_11_ANTENNA_DELAY_4 1
`define BEAM_11_ANTENNA_DELAY_5 10
`define BEAM_11_ANTENNA_DELAY_6 10
`define BEAM_11_ANTENNA_DELAY_7 9
`define BEAM_12_ANTENNA_DELAY_0 0
`define BEAM_12_ANTENNA_DELAY_1 11
`define BEAM_12_ANTENNA_DELAY_2 11
`define BEAM_12_ANTENNA_DELAY_3 10
`define BEAM_12_ANTENNA_DELAY_4 1
`define BEAM_12_ANTENNA_DELAY_5 11
`define BEAM_12_ANTENNA_DELAY_6 11
`define BEAM_12_ANTENNA_DELAY_7 10
`define BEAM_13_ANTENNA_DELAY_0 0
`define BEAM_13_ANTENNA_DELAY_1 12
`define BEAM_13_ANTENNA_DELAY_2 12
`define BEAM_13_ANTENNA_DELAY_3 12
`define BEAM_13_ANTENNA_DELAY_4 1
`define BEAM_13_ANTENNA_DELAY_5 12
`define BEAM_13_ANTENNA_DELAY_6 11
`define BEAM_13_ANTENNA_DELAY_7 11
`define BEAM_14_ANTENNA_DELAY_0 0
`define BEAM_14_ANTENNA_DELAY_1 12
`define BEAM_14_ANTENNA_DELAY_2 11
`define BEAM_14_ANTENNA_DELAY_3 11
`define BEAM_14_ANTENNA_DELAY_4 1
`define BEAM_14_ANTENNA_DELAY_5 12
`define BEAM_14_ANTENNA_DELAY_6 12
`define BEAM_14_ANTENNA_DELAY_7 12
`define BEAM_15_ANTENNA_DELAY_0 0
`define BEAM_15_ANTENNA_DELAY_1 13
`define BEAM_15_ANTENNA_DELAY_2 13
`define BEAM_15_ANTENNA_DELAY_3 13
`define BEAM_15_ANTENNA_DELAY_4 0
`define BEAM_15_ANTENNA_DELAY_5 13
`define BEAM_15_ANTENNA_DELAY_6 13
`define BEAM_15_ANTENNA_DELAY_7 13
`define BEAM_16_ANTENNA_DELAY_0 0
`define BEAM_16_ANTENNA_DELAY_1 14
`define BEAM_16_ANTENNA_DELAY_2 14
`define BEAM_16_ANTENNA_DELAY_3 14
`define BEAM_16_ANTENNA_DELAY_4 1
`define BEAM_16_ANTENNA_DELAY_5 15
`define BEAM_16_ANTENNA_DELAY_6 15
`define BEAM_16_ANTENNA_DELAY_7 15
`define BEAM_17_ANTENNA_DELAY_0 0
`define BEAM_17_ANTENNA_DELAY_1 15
`define BEAM_17_ANTENNA_DELAY_2 15
`define BEAM_17_ANTENNA_DELAY_3 15
`define BEAM_17_ANTENNA_DELAY_4 0
`define BEAM_17_ANTENNA_DELAY_5 14
`define BEAM_17_ANTENNA_DELAY_6 14
`define BEAM_17_ANTENNA_DELAY_7 14
`define BEAM_18_ANTENNA_DELAY_0 0
`define BEAM_18_ANTENNA_DELAY_1 15
`define BEAM_18_ANTENNA_DELAY_2 16
`define BEAM_18_ANTENNA_DELAY_3 17
`define BEAM_18_ANTENNA_DELAY_4 0
`define BEAM_18_ANTENNA_DELAY_5 15
`define BEAM_18_ANTENNA_DELAY_6 16
`define BEAM_18_ANTENNA_DELAY_7 17
`define BEAM_19_ANTENNA_DELAY_0 0
`define BEAM_19_ANTENNA_DELAY_1 16
`define BEAM_19_ANTENNA_DELAY_2 17
`define BEAM_19_ANTENNA_DELAY_3 18
`define BEAM_19_ANTENNA_DELAY_4 1
`define BEAM_19_ANTENNA_DELAY_5 17
`define BEAM_19_ANTENNA_DELAY_6 18
`define BEAM_19_ANTENNA_DELAY_7 18
`define BEAM_20_ANTENNA_DELAY_0 1
`define BEAM_20_ANTENNA_DELAY_1 17
`define BEAM_20_ANTENNA_DELAY_2 18
`define BEAM_20_ANTENNA_DELAY_3 18
`define BEAM_20_ANTENNA_DELAY_4 0
`define BEAM_20_ANTENNA_DELAY_5 16
`define BEAM_20_ANTENNA_DELAY_6 17
`define BEAM_20_ANTENNA_DELAY_7 18
`define BEAM_21_ANTENNA_DELAY_0 1
`define BEAM_21_ANTENNA_DELAY_1 17
`define BEAM_21_ANTENNA_DELAY_2 19
`define BEAM_21_ANTENNA_DELAY_3 20
`define BEAM_21_ANTENNA_DELAY_4 0
`define BEAM_21_ANTENNA_DELAY_5 17
`define BEAM_21_ANTENNA_DELAY_6 19
`define BEAM_21_ANTENNA_DELAY_7 20
`define BEAM_22_ANTENNA_DELAY_0 0
`define BEAM_22_ANTENNA_DELAY_1 17
`define BEAM_22_ANTENNA_DELAY_2 18
`define BEAM_22_ANTENNA_DELAY_3 20
`define BEAM_22_ANTENNA_DELAY_4 0
`define BEAM_22_ANTENNA_DELAY_5 18
`define BEAM_22_ANTENNA_DELAY_6 19
`define BEAM_22_ANTENNA_DELAY_7 21
`define BEAM_23_ANTENNA_DELAY_0 1
`define BEAM_23_ANTENNA_DELAY_1 19
`define BEAM_23_ANTENNA_DELAY_2 20
`define BEAM_23_ANTENNA_DELAY_3 22
`define BEAM_23_ANTENNA_DELAY_4 0
`define BEAM_23_ANTENNA_DELAY_5 18
`define BEAM_23_ANTENNA_DELAY_6 19
`define BEAM_23_ANTENNA_DELAY_7 21
`define BEAM_24_ANTENNA_DELAY_0 1
`define BEAM_24_ANTENNA_DELAY_1 20
`define BEAM_24_ANTENNA_DELAY_2 21
`define BEAM_24_ANTENNA_DELAY_3 23
`define BEAM_24_ANTENNA_DELAY_4 0
`define BEAM_24_ANTENNA_DELAY_5 20
`define BEAM_24_ANTENNA_DELAY_6 21
`define BEAM_24_ANTENNA_DELAY_7 23
`define BEAM_25_ANTENNA_DELAY_0 1
`define BEAM_25_ANTENNA_DELAY_1 21
`define BEAM_25_ANTENNA_DELAY_2 23
`define BEAM_25_ANTENNA_DELAY_3 25
`define BEAM_25_ANTENNA_DELAY_4 0
`define BEAM_25_ANTENNA_DELAY_5 20
`define BEAM_25_ANTENNA_DELAY_6 22
`define BEAM_25_ANTENNA_DELAY_7 24
`define BEAM_26_ANTENNA_DELAY_0 1
`define BEAM_26_ANTENNA_DELAY_1 20
`define BEAM_26_ANTENNA_DELAY_2 22
`define BEAM_26_ANTENNA_DELAY_3 24
`define BEAM_26_ANTENNA_DELAY_4 0
`define BEAM_26_ANTENNA_DELAY_5 21
`define BEAM_26_ANTENNA_DELAY_6 23
`define BEAM_26_ANTENNA_DELAY_7 25
`define BEAM_27_ANTENNA_DELAY_0 1
`define BEAM_27_ANTENNA_DELAY_1 22
`define BEAM_27_ANTENNA_DELAY_2 24
`define BEAM_27_ANTENNA_DELAY_3 26
`define BEAM_27_ANTENNA_DELAY_4 0
`define BEAM_27_ANTENNA_DELAY_5 22
`define BEAM_27_ANTENNA_DELAY_6 24
`define BEAM_27_ANTENNA_DELAY_7 26
`define BEAM_28_ANTENNA_DELAY_0 2
`define BEAM_28_ANTENNA_DELAY_1 23
`define BEAM_28_ANTENNA_DELAY_2 25
`define BEAM_28_ANTENNA_DELAY_3 28
`define BEAM_28_ANTENNA_DELAY_4 0
`define BEAM_28_ANTENNA_DELAY_5 22
`define BEAM_28_ANTENNA_DELAY_6 25
`define BEAM_28_ANTENNA_DELAY_7 27
`define BEAM_29_ANTENNA_DELAY_0 1
`define BEAM_29_ANTENNA_DELAY_1 22
`define BEAM_29_ANTENNA_DELAY_2 25
`define BEAM_29_ANTENNA_DELAY_3 27
`define BEAM_29_ANTENNA_DELAY_4 0
`define BEAM_29_ANTENNA_DELAY_5 23
`define BEAM_29_ANTENNA_DELAY_6 25
`define BEAM_29_ANTENNA_DELAY_7 28
`define BEAM_30_ANTENNA_DELAY_0 2
`define BEAM_30_ANTENNA_DELAY_1 24
`define BEAM_30_ANTENNA_DELAY_2 26
`define BEAM_30_ANTENNA_DELAY_3 29
`define BEAM_30_ANTENNA_DELAY_4 0
`define BEAM_30_ANTENNA_DELAY_5 24
`define BEAM_30_ANTENNA_DELAY_6 26
`define BEAM_30_ANTENNA_DELAY_7 29
`define BEAM_31_ANTENNA_DELAY_0 2
`define BEAM_31_ANTENNA_DELAY_1 25
`define BEAM_31_ANTENNA_DELAY_2 28
`define BEAM_31_ANTENNA_DELAY_3 31
`define BEAM_31_ANTENNA_DELAY_4 0
`define BEAM_31_ANTENNA_DELAY_5 24
`define BEAM_31_ANTENNA_DELAY_6 27
`define BEAM_31_ANTENNA_DELAY_7 30
`define BEAM_32_ANTENNA_DELAY_0 2
`define BEAM_32_ANTENNA_DELAY_1 24
`define BEAM_32_ANTENNA_DELAY_2 27
`define BEAM_32_ANTENNA_DELAY_3 30
`define BEAM_32_ANTENNA_DELAY_4 0
`define BEAM_32_ANTENNA_DELAY_5 25
`define BEAM_32_ANTENNA_DELAY_6 28
`define BEAM_32_ANTENNA_DELAY_7 31
`define BEAM_33_ANTENNA_DELAY_0 2
`define BEAM_33_ANTENNA_DELAY_1 26
`define BEAM_33_ANTENNA_DELAY_2 29
`define BEAM_33_ANTENNA_DELAY_3 32
`define BEAM_33_ANTENNA_DELAY_4 0
`define BEAM_33_ANTENNA_DELAY_5 26
`define BEAM_33_ANTENNA_DELAY_6 29
`define BEAM_33_ANTENNA_DELAY_7 32
`define BEAM_34_ANTENNA_DELAY_0 2
`define BEAM_34_ANTENNA_DELAY_1 27
`define BEAM_34_ANTENNA_DELAY_2 31
`define BEAM_34_ANTENNA_DELAY_3 34
`define BEAM_34_ANTENNA_DELAY_4 0
`define BEAM_34_ANTENNA_DELAY_5 27
`define BEAM_34_ANTENNA_DELAY_6 30
`define BEAM_34_ANTENNA_DELAY_7 33
`define BEAM_35_ANTENNA_DELAY_0 2
`define BEAM_35_ANTENNA_DELAY_1 27
`define BEAM_35_ANTENNA_DELAY_2 30
`define BEAM_35_ANTENNA_DELAY_3 33
`define BEAM_35_ANTENNA_DELAY_4 0
`define BEAM_35_ANTENNA_DELAY_5 27
`define BEAM_35_ANTENNA_DELAY_6 31
`define BEAM_35_ANTENNA_DELAY_7 34
`define BEAM_36_ANTENNA_DELAY_0 2
`define BEAM_36_ANTENNA_DELAY_1 28
`define BEAM_36_ANTENNA_DELAY_2 32
`define BEAM_36_ANTENNA_DELAY_3 35
`define BEAM_36_ANTENNA_DELAY_4 0
`define BEAM_36_ANTENNA_DELAY_5 28
`define BEAM_36_ANTENNA_DELAY_6 32
`define BEAM_36_ANTENNA_DELAY_7 35
`define BEAM_37_ANTENNA_DELAY_0 3
`define BEAM_37_ANTENNA_DELAY_1 29
`define BEAM_37_ANTENNA_DELAY_2 33
`define BEAM_37_ANTENNA_DELAY_3 37
`define BEAM_37_ANTENNA_DELAY_4 0
`define BEAM_37_ANTENNA_DELAY_5 29
`define BEAM_37_ANTENNA_DELAY_6 33
`define BEAM_37_ANTENNA_DELAY_7 36
`define BEAM_38_ANTENNA_DELAY_0 2
`define BEAM_38_ANTENNA_DELAY_1 29
`define BEAM_38_ANTENNA_DELAY_2 33
`define BEAM_38_ANTENNA_DELAY_3 36
`define BEAM_38_ANTENNA_DELAY_4 0
`define BEAM_38_ANTENNA_DELAY_5 29
`define BEAM_38_ANTENNA_DELAY_6 33
`define BEAM_38_ANTENNA_DELAY_7 37
`define BEAM_39_ANTENNA_DELAY_0 3
`define BEAM_39_ANTENNA_DELAY_1 30
`define BEAM_39_ANTENNA_DELAY_2 34
`define BEAM_39_ANTENNA_DELAY_3 38
`define BEAM_39_ANTENNA_DELAY_4 0
`define BEAM_39_ANTENNA_DELAY_5 30
`define BEAM_39_ANTENNA_DELAY_6 34
`define BEAM_39_ANTENNA_DELAY_7 38
`define BEAM_40_ANTENNA_DELAY_0 3
`define BEAM_40_ANTENNA_DELAY_1 31
`define BEAM_40_ANTENNA_DELAY_2 36
`define BEAM_40_ANTENNA_DELAY_3 40
`define BEAM_40_ANTENNA_DELAY_4 0
`define BEAM_40_ANTENNA_DELAY_5 31
`define BEAM_40_ANTENNA_DELAY_6 35
`define BEAM_40_ANTENNA_DELAY_7 40
`define BEAM_41_ANTENNA_DELAY_0 3
`define BEAM_41_ANTENNA_DELAY_1 31
`define BEAM_41_ANTENNA_DELAY_2 35
`define BEAM_41_ANTENNA_DELAY_3 40
`define BEAM_41_ANTENNA_DELAY_4 0
`define BEAM_41_ANTENNA_DELAY_5 31
`define BEAM_41_ANTENNA_DELAY_6 36
`define BEAM_41_ANTENNA_DELAY_7 40
`define BEAM_42_ANTENNA_DELAY_0 3
`define BEAM_42_ANTENNA_DELAY_1 32
`define BEAM_42_ANTENNA_DELAY_2 37
`define BEAM_42_ANTENNA_DELAY_3 41
`define BEAM_42_ANTENNA_DELAY_4 0
`define BEAM_42_ANTENNA_DELAY_5 32
`define BEAM_42_ANTENNA_DELAY_6 37
`define BEAM_42_ANTENNA_DELAY_7 41
`define BEAM_43_ANTENNA_DELAY_0 4
`define BEAM_43_ANTENNA_DELAY_1 33
`define BEAM_43_ANTENNA_DELAY_2 38
`define BEAM_43_ANTENNA_DELAY_3 43
`define BEAM_43_ANTENNA_DELAY_4 0
`define BEAM_43_ANTENNA_DELAY_5 33
`define BEAM_43_ANTENNA_DELAY_6 38
`define BEAM_43_ANTENNA_DELAY_7 43
`define BEAM_44_ANTENNA_DELAY_0 3
`define BEAM_44_ANTENNA_DELAY_1 33
`define BEAM_44_ANTENNA_DELAY_2 38
`define BEAM_44_ANTENNA_DELAY_3 43
`define BEAM_44_ANTENNA_DELAY_4 0
`define BEAM_44_ANTENNA_DELAY_5 34
`define BEAM_44_ANTENNA_DELAY_6 38
`define BEAM_44_ANTENNA_DELAY_7 43
`define BEAM_45_ANTENNA_DELAY_0 4
`define BEAM_45_ANTENNA_DELAY_1 34
`define BEAM_45_ANTENNA_DELAY_2 39
`define BEAM_45_ANTENNA_DELAY_3 45
`define BEAM_45_ANTENNA_DELAY_4 0
`define BEAM_45_ANTENNA_DELAY_5 34
`define BEAM_45_ANTENNA_DELAY_6 39
`define BEAM_45_ANTENNA_DELAY_7 45
`define MAX_ANTENNA_DELAY_0 4
`define MAX_ANTENNA_DELAY_4 3
