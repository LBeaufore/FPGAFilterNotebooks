`define BEAM_0_ANTENNA_DELAYS { 1 4 2 0 3 4 2 0 }
`define BEAM_1_ANTENNA_DELAYS { 0 5 3 1 2 4 2 0 }
`define BEAM_2_ANTENNA_DELAYS { 0 4 2 0 2 5 3 1 }
`define BEAM_3_ANTENNA_DELAYS { 0 5 4 2 2 5 4 2 }
`define BEAM_4_ANTENNA_DELAYS { 0 7 5 4 2 6 5 3 }
`define BEAM_5_ANTENNA_DELAYS { 0 6 5 3 2 7 5 4 }
`define BEAM_6_ANTENNA_DELAYS { 0 8 6 5 2 8 6 5 }
`define BEAM_7_ANTENNA_DELAYS { 0 8 7 6 1 7 6 5 }
`define BEAM_8_ANTENNA_DELAYS { 0 8 7 6 2 9 8 7 }
`define BEAM_9_ANTENNA_DELAYS { 0 10 9 8 2 10 9 8 }
`define BEAM_10_ANTENNA_DELAYS { 0 10 10 9 1 9 9 8 }
`define BEAM_12_ANTENNA_DELAYS { 0 11 11 10 1 11 11 10 }
`define BEAM_13_ANTENNA_DELAYS { 0 12 12 12 1 12 11 11 }
`define BEAM_14_ANTENNA_DELAYS { 0 12 11 11 1 12 12 12 }
`define BEAM_15_ANTENNA_DELAYS { 0 13 13 13 0 13 13 13 }
`define BEAM_16_ANTENNA_DELAYS { 0 14 14 14 1 15 15 15 }
`define BEAM_17_ANTENNA_DELAYS { 0 15 15 15 0 14 14 14 }
`define BEAM_18_ANTENNA_DELAYS { 0 15 16 17 0 15 16 17 }
`define BEAM_19_ANTENNA_DELAYS { 0 16 17 18 1 17 18 18 }
`define BEAM_20_ANTENNA_DELAYS { 1 17 18 18 0 16 17 18 }
`define BEAM_21_ANTENNA_DELAYS { 1 17 19 20 0 17 19 20 }
`define BEAM_22_ANTENNA_DELAYS { 0 17 18 20 0 18 19 21 }
`define BEAM_23_ANTENNA_DELAYS { 1 19 20 22 0 18 19 21 }
`define BEAM_24_ANTENNA_DELAYS { 1 20 21 23 0 20 21 23 }
`define BEAM_25_ANTENNA_DELAYS { 1 21 23 25 0 20 22 24 }
`define BEAM_26_ANTENNA_DELAYS { 1 20 22 24 0 21 23 25 }
`define BEAM_27_ANTENNA_DELAYS { 1 22 24 26 0 22 24 26 }
`define BEAM_28_ANTENNA_DELAYS { 2 23 25 28 0 22 25 27 }
`define BEAM_29_ANTENNA_DELAYS { 1 22 25 27 0 23 25 28 }
`define BEAM_30_ANTENNA_DELAYS { 2 24 26 29 0 24 26 29 }
`define BEAM_31_ANTENNA_DELAYS { 2 25 28 31 0 24 27 30 }
`define BEAM_32_ANTENNA_DELAYS { 2 24 27 30 0 25 28 31 }
`define BEAM_33_ANTENNA_DELAYS { 2 26 29 32 0 26 29 32 }
`define BEAM_34_ANTENNA_DELAYS { 2 27 31 34 0 27 30 33 }
`define BEAM_35_ANTENNA_DELAYS { 2 27 30 33 0 27 31 34 }
`define BEAM_36_ANTENNA_DELAYS { 2 28 32 35 0 28 32 35 }
`define BEAM_37_ANTENNA_DELAYS { 3 29 33 37 0 29 33 36 }
`define BEAM_38_ANTENNA_DELAYS { 2 29 33 36 0 29 33 37 }
`define BEAM_39_ANTENNA_DELAYS { 3 30 34 38 0 30 34 38 }
`define BEAM_40_ANTENNA_DELAYS { 3 31 36 40 0 31 35 40 }
`define BEAM_41_ANTENNA_DELAYS { 3 31 35 40 0 31 36 40 }
`define BEAM_42_ANTENNA_DELAYS { 3 32 37 41 0 32 37 41 }
`define BEAM_43_ANTENNA_DELAYS { 4 33 38 43 0 33 38 43 }
`define BEAM_44_ANTENNA_DELAYS { 3 33 38 43 0 34 38 43 }
`define BEAM_45_ANTENNA_DELAYS { 4 34 39 45 0 34 39 45 }
`define MAX_ANTENNA_DELAY_0 4
`define MAX_ANTENNA_DELAY_1 34
`define MAX_ANTENNA_DELAY_2 39
`define MAX_ANTENNA_DELAY_3 45
`define MAX_ANTENNA_DELAY_4 3
`define MAX_ANTENNA_DELAY_5 34
`define MAX_ANTENNA_DELAY_6 39
`define MAX_ANTENNA_DELAY_7 45
